./tests.verify: test performed on 2004.03.14 


#### Test: ./tests.verify running commontasks.py 
Hello Pipe World
./commontasks.py : cannot read file 'qqq'
An exception of type
  exceptions.IOError 
occurred, with value
   [Errno 2] No such file or directory: 'qqq'
arglist= ['myarg1', 'displacement', 'tmp.ps']
filename= myarg1  plottitle= displacement  psfile= tmp.ps
arglist= ['myarg1', 'displacement', 'tmp.ps', 'myvar2']
entry is  myarg1
entry is  displacement
entry is  tmp.ps
entry is  myvar2
In-place manipulation of array entries:
A[0]=1.2
A[1]=-3.4
A[2]=5.5
A[3]=-9
A[4]=100
No negative numbers:
A[0]=1.2
A[1]=0
A[2]=5.5
A[3]=0
A[4]=100
a 'foreach'-type loop does not work:
A[0]=1.2
A[1]=-3.4
A[2]=5.5
A[3]=-9
A[4]=100

split with re.split:
words1[0] = "iteration"
words1[1] = "12:"
words1[2] = "eps="
words1[3] = "1.245E-05"

split with string.split instead:
words1[0] = "iteration"
words1[2] = "12:"
words1[4] = "eps="
words1[6] = "1.245E-05"
newline1 is now [ iteration#12:#eps=#1.245E-05 ]
words2[0]=.myc_12
words2[1]=displacement
words2[2]=u(x,3.1415)
words2[3]=  no upwinding
['white', 'space', 'of', 'varying', 'length']
['white', 'space', '', '', 'of', 'varying', '', '', '', 'length']
Yes, matched regex= <_sre.SRE_Match object at 0x4022eaa0>
regex sub:
#!/usr/bin/env python
import sys, math       # load system and math module
r = float(sys.argv[1]) # extract the 1st command-line arg.
s = math.sin(r)
print "Hello, World! sin(" + str(r) + ")=" + str(s)



Testing dictionaries:

len(myargs)= 6
The option --myopt is not registered
The option -9.9 is not registered
dictionary: cmlargs, key= -tstop  value= 6.1
dictionary: cmlargs, key= -c_in_H  value= 9.8
cmlargs['-c_in_H']=9.8
cmlargs['-tstop']=6.1




Python lacks auto convert of strings-numbers
a =  0.6
hw.py is a plain file
stat:  33261
stat:  68938
stat:  778
stat:  1
stat:  8029
stat:  8029
stat:  202
stat:  1079261774
stat:  1071617117
stat:  1073569782
hw.py is a regular file with 202 bytes and last accessed 1079261774
0.16Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1571.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2180.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1614.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/solaris_thr.gif
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2204.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2215.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2219.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1639.xbm
0.04Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2230.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/thread_stack.gif
0.05Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2282.xbm
0.04Mb /work/scripting/doc/c/tutorial/C/node1.html
0.02Mb /work/scripting/doc/c/tutorial/C/node2.html
0.02Mb /work/scripting/doc/c/tutorial/C/node3.html
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing51.xbm
0.04Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing54.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing58.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/node4.html
0.01Mb /work/scripting/doc/c/tutorial/C/node6.html
0.12Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2355.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node8.html
0.01Mb /work/scripting/doc/c/tutorial/C/node9.html
0.01Mb /work/scripting/doc/c/tutorial/C/subsection2_19_3_2.html
0.01Mb /work/scripting/doc/c/tutorial/C/notes.gif
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2388.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing162.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing170.xbm
0.06Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2412.xbm
0.06Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2416.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1830.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing224.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing234.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing245.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/node10.html
0.02Mb /work/scripting/doc/c/tutorial/C/mthread.gif
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing277.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing279.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node11.html
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1237.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1930.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node12.html
0.01Mb /work/scripting/doc/c/tutorial/C/node13.html
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1948.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node14.html
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1958.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node16.html
0.02Mb /work/scripting/doc/c/tutorial/C/node18.html
0.04Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing344.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node19.html
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing351.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing353.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/node20.html
0.01Mb /work/scripting/doc/c/tutorial/C/node22.html
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing398.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/node24.html
0.04Mb /work/scripting/doc/c/tutorial/C/node25.html
0.05Mb /work/scripting/doc/c/tutorial/C/CE.html
0.04Mb /work/scripting/doc/c/tutorial/C/node26.html
0.01Mb /work/scripting/doc/c/tutorial/C/CDE.gif
0.04Mb /work/scripting/doc/c/tutorial/C/node27.html
0.03Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing431.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Courseware.txt
0.08Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Develop.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Tutor.txt
0.05Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Design.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Stats.txt
0.05Mb /work/scripting/doc/c/tutorial/C/CEILIDH/ASQA.txt
0.01Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Qu-ans.txt
0.03Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Student.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes1.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes2.txt
0.01Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes3.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes4.txt
0.03Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes5.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes6.txt
0.03Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes7.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/notes8.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Overview.txt
0.03Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Install.txt
0.02Mb /work/scripting/doc/c/tutorial/C/CEILIDH/Teacher.txt
0.02Mb /work/scripting/doc/c/tutorial/C/node28.html
0.07Mb /work/scripting/doc/c/tutorial/C/node29.html
0.03Mb /work/scripting/doc/c/tutorial/C/node30.html
0.05Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing471.xbm
0.05Mb /work/scripting/doc/c/tutorial/C/node31.html
0.12Mb /work/scripting/doc/c/tutorial/C/node32.html
0.04Mb /work/scripting/doc/c/tutorial/C/node33.html
0.05Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1455.xbm
0.04Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2050.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/node34.html
0.02Mb /work/scripting/doc/c/tutorial/C/node35.html
0.01Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1475.xbm
0.18Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2074.xbm
0.03Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2077.xbm
0.08Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing2091.xbm
0.01Mb /work/scripting/doc/c/tutorial/C/mainw.gif
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1501.xbm
0.04Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1522.xbm
0.02Mb /work/scripting/doc/c/tutorial/C/_17661_tabbing1532.xbm
0.02Mb /work/scripting/doc/tk/font.html
0.03Mb /work/scripting/doc/tk/options.html
0.04Mb /work/scripting/doc/tk/menu.html
0.02Mb /work/scripting/doc/tk/winfo.html
0.02Mb /work/scripting/doc/tk/scrollbar.html
0.01Mb /work/scripting/doc/tk/menubutton.html
0.03Mb /work/scripting/doc/tk/listbox.html
0.01Mb /work/scripting/doc/tk/button.html
0.02Mb /work/scripting/doc/tk/photo.html
0.02Mb /work/scripting/doc/tk/grid.html
0.09Mb /work/scripting/doc/tk/text.html
0.02Mb /work/scripting/doc/tk/scale.html
0.01Mb /work/scripting/doc/tk/place.html
0.01Mb /work/scripting/doc/tk/toplevel.html
0.01Mb /work/scripting/doc/tk/pack.html
0.09Mb /work/scripting/doc/tk/canvas.html
0.02Mb /work/scripting/doc/tk/radiobutton.html
0.01Mb /work/scripting/doc/tk/message.html
0.03Mb /work/scripting/doc/tk/wm.html
0.02Mb /work/scripting/doc/tk/event.html
0.03Mb /work/scripting/doc/tk/entry.html
0.02Mb /work/scripting/doc/tk/bind.html
0.02Mb /work/scripting/doc/tk/checkbutton.html
0.41Mb /work/scripting/doc/f77/F77-programming.html
0.01Mb /work/scripting/doc/cvs/cvs_toc.html
0.02Mb /work/scripting/doc/cvs/cvsintro.html
0.03Mb /work/scripting/doc/cvs/cvs_10.html
0.01Mb /work/scripting/doc/cvs/cvs_12.html
0.10Mb /work/scripting/doc/cvs/cvs_16.html
0.03Mb /work/scripting/doc/cvs/cvs_17.html
0.04Mb /work/scripting/doc/cvs/cvs_18.html
0.02Mb /work/scripting/doc/cvs/cvs_21.html
0.02Mb /work/scripting/doc/cvs/cvs_1.html
0.03Mb /work/scripting/doc/cvs/cvs_index.html
0.07Mb /work/scripting/doc/cvs/cvs_2.html
0.01Mb /work/scripting/doc/cvs/cvs_4.html
0.02Mb /work/scripting/doc/cvs/cvs_5.html
0.02Mb /work/scripting/doc/cvs/cvs_7.html
0.08Mb /work/scripting/doc/etc/mpeg_encode_userguide.ps
0.11Mb /work/scripting/doc/perl/perl5-quickref.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perltie.html
0.07Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq4.html
0.06Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq5.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq6.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq7.html
0.03Mb /work/scripting/doc/perl/Perl-FAQ/perlhist.html
0.06Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq8.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq9.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlxstut.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perllol.html
0.06Mb /work/scripting/doc/perl/Perl-FAQ/perlsub.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perlvar.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlbot.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlref.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perlmodlib.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlform.html
0.08Mb /work/scripting/doc/perl/Perl-FAQ/perlcall.html
0.07Mb /work/scripting/doc/perl/Perl-FAQ/perlipc.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perlembed.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlpod.html
0.09Mb /work/scripting/doc/perl/Perl-FAQ/perlop.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq.html
0.03Mb /work/scripting/doc/perl/Perl-FAQ/perlmod.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlrun.html
0.06Mb /work/scripting/doc/perl/Perl-FAQ/perldelta.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perltrap.html
0.05Mb /work/scripting/doc/perl/Perl-FAQ/perlre.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perldsc.html
0.03Mb /work/scripting/doc/perl/Perl-FAQ/perlsec.html
0.07Mb /work/scripting/doc/perl/Perl-FAQ/perlxs.html
0.23Mb /work/scripting/doc/perl/Perl-FAQ/perltoc.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlsyn.html
0.06Mb /work/scripting/doc/perl/Perl-FAQ/perllocale.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlstyle.html
0.17Mb /work/scripting/doc/perl/Perl-FAQ/perlguts.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perldata.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getgrgid.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getnetbyname.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getprotoent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endhostent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/sort.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/defined.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getservbyport.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getgrnam.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getprotobynumber.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/sethostent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endservent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getnetbyaddr.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endprotoent.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/index.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getpwnam.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/exec.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/open.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/split.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endnetent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/setservent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/setprotoent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/sprintf.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/gethostbyname.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/flock.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/gethostent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getservbyname.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endgrent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getpwuid.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/setgrent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getprotobyname.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/setnetent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/use.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/pack.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/eval.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getgrent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/endpwent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getservent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/gethostbyaddr.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/setpwent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getpwent.html
0.01Mb /work/scripting/doc/perl/Perl-FAQ/perlfunc/getnetent.html
0.08Mb /work/scripting/doc/perl/Perl-FAQ/perldebug.html
0.09Mb /work/scripting/doc/perl/Perl-FAQ/perltoot.html
0.02Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq1.html
0.03Mb /work/scripting/doc/perl/Perl-FAQ/perlobj.html
0.03Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq2.html
0.16Mb /work/scripting/doc/perl/Perl-FAQ/perldiag.html
0.04Mb /work/scripting/doc/perl/Perl-FAQ/perlfaq3.html
0.01Mb /work/scripting/doc/swig/manual/Arguments.html
0.04Mb /work/scripting/doc/swig/manual/Library.html
0.10Mb /work/scripting/doc/swig/manual/SWIGPlus.html
0.02Mb /work/scripting/doc/swig/manual/Advanced.html
0.08Mb /work/scripting/doc/swig/manual/Typemaps.html
0.09Mb /work/scripting/doc/swig/manual/Extending.html
0.13Mb /work/scripting/doc/swig/manual/Java.html
0.07Mb /work/scripting/doc/swig/manual/Perl5.html
0.02Mb /work/scripting/doc/swig/manual/Guile.html
0.08Mb /work/scripting/doc/swig/manual/Tcl.html
0.08Mb /work/scripting/doc/swig/manual/Ruby.html
0.03Mb /work/scripting/doc/swig/manual/Varargs.html
0.01Mb /work/scripting/doc/swig/manual/Introduction.html
0.02Mb /work/scripting/doc/swig/manual/Ocaml.html
0.08Mb /work/scripting/doc/swig/manual/SWIG.html
0.02Mb /work/scripting/doc/swig/manual/Customization.html
0.01Mb /work/scripting/doc/swig/manual/Warnings.html
0.09Mb /work/scripting/doc/swig/manual/Python.html
0.02Mb /work/scripting/doc/swig/manual/Php.html
0.04Mb /work/scripting/doc/swig/manual/Contents.html
0.01Mb /work/scripting/doc/swig/manual/Scripting.html
0.40Mb /work/scripting/doc/unix/unix_intro.html
0.04Mb /work/scripting/doc/latex/intro/textcomp.ps
0.02Mb /work/scripting/doc/latex/intro/reports.html
0.02Mb /work/scripting/doc/latex/intro/LaTeX_intro.html
0.01Mb /work/scripting/doc/latex/intro/teTeX/help/faq/uktug-faq/index.html
0.07Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctd.html
0.10Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cte.html
0.08Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctf.html
0.05Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctg.html
0.04Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cth.html
0.03Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cti.html
0.01Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctj.html
0.02Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctk.html
0.10Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctl.html
0.04Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctn.html
0.03Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cto.html
0.11Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctp.html
0.01Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctq.html
0.05Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctr.html
0.10Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cts.html
0.30Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctbrief.html
0.13Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctt.html
0.04Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctu.html
0.02Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctv.html
0.04Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctw.html
0.02Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctx.html
0.02Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cty.html
0.12Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctfull.html.gz
0.05Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctindex.html
0.19Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cthier.html
1.39Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctfull.html
0.12Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/cta.html
0.07Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctb.html
0.13Mb /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctc.html
2.82Mb /work/scripting/doc/latex/intro/teTeX/context/base/ms-cb-en.pdf
0.32Mb /work/scripting/doc/latex/intro/teTeX/context/base/setup-en.pdf
0.39Mb /work/scripting/doc/latex/intro/teTeX/metapost/base/mpgraph.ps
0.79Mb /work/scripting/doc/latex/intro/teTeX/metapost/base/mpman.ps
0.02Mb /work/scripting/doc/latex/intro/teTeX/fonts/ae/COPYING
0.01Mb /work/scripting/doc/latex/intro/teTeX/fonts/ec/changelog
0.01Mb /work/scripting/doc/latex/intro/teTeX/fonts/pl/readme.eng
0.01Mb /work/scripting/doc/latex/intro/teTeX/fonts/pl/readme.pol
0.02Mb /work/scripting/doc/latex/intro/teTeX/fonts/fontname/ChangeLog
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/base/manual.err
0.10Mb /work/scripting/doc/latex/intro/teTeX/latex/base/compan.err
0.08Mb /work/scripting/doc/latex/intro/teTeX/latex/base/begleit.err
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/base/manifest.txt
0.23Mb /work/scripting/doc/latex/intro/teTeX/latex/base/changes.txt
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/latex2e-html/ltx-2.html
0.08Mb /work/scripting/doc/latex/intro/teTeX/latex/amslatex/testmath.tex
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/amslatex/amslatex.bug
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/amslatex/diff12.tex
0.05Mb /work/scripting/doc/latex/intro/teTeX/latex/amslatex/instr-l.tex
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/amslatex/technote.tex
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/custom-bib/shorthnd.tex
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/custom-bib/geophys.tex
0.32Mb /work/scripting/doc/latex/intro/teTeX/latex/graphics/grfguide.ps
2.31Mb /work/scripting/doc/latex/intro/teTeX/latex/graphics/epslatex.ps
0.03Mb /work/scripting/doc/latex/intro/teTeX/latex/tools/changes.txt
0.43Mb /work/scripting/doc/latex/intro/teTeX/latex/fancyvrb/fancyvrb.ps
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/seminar/sem-read.me
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/seminar/semsamp2.tex
0.03Mb /work/scripting/doc/latex/intro/teTeX/latex/seminar/Seminar-Bugs.html
0.06Mb /work/scripting/doc/latex/intro/teTeX/latex/seminar/Seminar-FAQ.html
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/minitoc/minitoc-ex.tex
0.15Mb /work/scripting/doc/latex/intro/teTeX/latex/general/guide.ps
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/mathtime/test11p.tex
0.31Mb /work/scripting/doc/latex/intro/teTeX/latex/carlisle/colortbl.ps
0.33Mb /work/scripting/doc/latex/intro/teTeX/latex/rotating/examples.ps
0.01Mb /work/scripting/doc/latex/intro/teTeX/latex/rotating/examples.tex
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/rotating/cat.eps
0.08Mb /work/scripting/doc/latex/intro/teTeX/latex/rotfloat/examples.ps
0.29Mb /work/scripting/doc/latex/intro/teTeX/latex/psfrag/pfgguide.ps
0.33Mb /work/scripting/doc/latex/intro/teTeX/latex/oberdiek/hypbmsec.pdf
0.29Mb /work/scripting/doc/latex/intro/teTeX/latex/oberdiek/twoopt.pdf
0.37Mb /work/scripting/doc/latex/intro/teTeX/latex/oberdiek/alphalph.pdf
0.34Mb /work/scripting/doc/latex/intro/teTeX/latex/oberdiek/pagesel.pdf
0.05Mb /work/scripting/doc/latex/intro/teTeX/latex/styles/index.doc
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/styles/readme.fp
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/floatflt/floatexm.tex
0.18Mb /work/scripting/doc/latex/intro/teTeX/latex/hyperref/manual.pdf
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/mdwtools/README
0.02Mb /work/scripting/doc/latex/intro/teTeX/latex/mdwtools/COPYING
0.03Mb /work/scripting/doc/latex/intro/teTeX/tetex/teTeX-FAQ
0.04Mb /work/scripting/doc/latex/intro/teTeX/index.html
0.01Mb /work/scripting/doc/latex/intro/teTeX/amstex/joyerr.tex
0.98Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/doc-fill.ps
0.01Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/CHANGES
0.12Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/pst-usr1.ps
0.13Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/pst-usr2.ps
0.15Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/pst-usr3.ps
0.11Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/pst-usr4.ps
0.19Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/betadoc1.ps
0.24Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/betadoc2.ps
0.06Mb /work/scripting/doc/latex/intro/teTeX/generic/pstricks/obsolete/pst-quik.ps
0.06Mb /work/scripting/doc/latex/intro/teTeX/generic/babel/changes.txt
0.67Mb /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyguide.ps
1.86Mb /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyrefer.ps
0.02Mb /work/scripting/doc/latex/intro/teTeX/generic/xypic/COPYING
0.01Mb /work/scripting/doc/latex/intro/teTeX/generic/texdraw/txdexamp.latex
0.43Mb /work/scripting/doc/latex/intro/teTeX/generic/texdraw/texdraw.ps
0.25Mb /work/scripting/doc/latex/intro/teTeX/pdftex/base/pdftexman.pdf
0.09Mb /work/scripting/doc/latex/intro/teTeX/pdftex/base/pdfTeX-FAQ.pdf
0.04Mb /work/scripting/doc/latex/intro/teTeX/newhelpindex.html
0.17Mb /work/scripting/doc/latex/intro/symbols.ps
0.20Mb /work/scripting/doc/latex/intro/psfrag.ps
1.01Mb /work/scripting/doc/latex/intro/ltxprimer-1.0.pdf
0.06Mb /work/scripting/doc/latex/intro/quickrep.pdf
0.25Mb /work/scripting/doc/latex/intro/lablet98man.ps
0.03Mb /work/scripting/doc/latex/intro/fonts.html
1.31Mb /work/scripting/doc/latex/intro/tipaman.pdf
0.02Mb /work/scripting/doc/latex/intro/index.html
0.17Mb /work/scripting/doc/latex/intro/colortbl.ps
0.02Mb /work/scripting/doc/latex/intro/latex2html/node47.html
0.02Mb /work/scripting/doc/latex/intro/latex2html/node6.html
0.03Mb /work/scripting/doc/latex/intro/latex2html/img8.gif
0.01Mb /work/scripting/doc/latex/intro/latex2html/node34.html
0.01Mb /work/scripting/doc/latex/intro/latex2html/node36.html
0.01Mb /work/scripting/doc/latex/intro/latex2html/node41.html
0.46Mb /work/scripting/doc/latex/intro/prosper-doc.pdf
0.11Mb /work/scripting/doc/latex/intro/contour.ps
0.10Mb /work/scripting/doc/latex/intro/prosper-tour.pdf
0.01Mb /work/scripting/doc/latex/intro/extending_latex.html
0.24Mb /work/scripting/doc/latex/intro/rotating.ps
0.02Mb /work/scripting/doc/latex/intro/makingWWWdocs.html
0.02Mb /work/scripting/doc/latex/intro/latex_maths+pix/node6.html
0.77Mb /work/scripting/doc/latex/intro/epslatex.ps
0.03Mb /work/scripting/doc/latex/intro/latex_advanced/node14.html
0.04Mb /work/scripting/doc/ImageMagick/www/api/image.html
0.02Mb /work/scripting/doc/ImageMagick/www/api/types/Enumerations.html
0.01Mb /work/scripting/doc/ImageMagick/www/api/types/ImageInfo.html
0.02Mb /work/scripting/doc/ImageMagick/www/api/types/Image.html
0.01Mb /work/scripting/doc/ImageMagick/www/api/mac.html
0.02Mb /work/scripting/doc/ImageMagick/www/api/widget.html
0.02Mb /work/scripting/doc/ImageMagick/www/api/utility.html
0.06Mb /work/scripting/doc/ImageMagick/www/api/xwindows.html
0.03Mb /work/scripting/doc/ImageMagick/www/api/effects.html
0.02Mb /work/scripting/doc/ImageMagick/www/api/blob.html
0.01Mb /work/scripting/doc/ImageMagick/www/api/compress.html
0.02Mb /work/scripting/doc/ImageMagick/www/miff.html
0.03Mb /work/scripting/doc/ImageMagick/www/Magick.html
0.05Mb /work/scripting/doc/ImageMagick/www/perl.html
0.05Mb /work/scripting/doc/ImageMagick/www/install.html
0.02Mb /work/scripting/doc/ImageMagick/www/quantize.html
0.06Mb /work/scripting/doc/ImageMagick/www/montage.html
0.07Mb /work/scripting/doc/ImageMagick/www/mogrify.html
0.04Mb /work/scripting/doc/ImageMagick/www/combine.html
0.04Mb /work/scripting/doc/ImageMagick/www/import.html
0.08Mb /work/scripting/doc/ImageMagick/www/convert.html
0.02Mb /work/scripting/doc/ImageMagick/www/formats.html
0.02Mb /work/scripting/doc/ImageMagick/www/xtp.html
0.05Mb /work/scripting/doc/ImageMagick/www/Changelog.html
0.04Mb /work/scripting/doc/ImageMagick/www/animate.html
0.13Mb /work/scripting/doc/ImageMagick/www/display.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/fig/sample9.6a.png
0.02Mb /work/scripting/doc/gnuplot/Kawano/fig/sample9.6b.png
0.02Mb /work/scripting/doc/gnuplot/Kawano/fig/sample8.3d.jpg
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/index.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/besj0.eps
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/besj1.eps
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/index-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/besy0.eps
0.01Mb /work/scripting/doc/gnuplot/Kawano/esub/besy1.eps
0.03Mb /work/scripting/doc/gnuplot/Kawano/esub/figure1.ps
0.03Mb /work/scripting/doc/gnuplot/Kawano/esub/figure2.ps
0.03Mb /work/scripting/doc/gnuplot/Kawano/esub/figure3.ps
0.03Mb /work/scripting/doc/gnuplot/Kawano/esub/figure4.ps
0.08Mb /work/scripting/doc/gnuplot/Kawano/esub/figure5.ps
0.03Mb /work/scripting/doc/gnuplot/Kawano/esub/figure6.ps
0.01Mb /work/scripting/doc/gnuplot/Kawano/set-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot3d-e.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/datafile2.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/datafile.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/postscript.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/image/world.png
0.07Mb /work/scripting/doc/gnuplot/Kawano/image/graph-new.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/style-e.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/intro/plotexp.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/intro/manyfigure.png
0.02Mb /work/scripting/doc/gnuplot/Kawano/intro/basic-e.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/intro/basic.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/working.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/working-e.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/intro/plotexp-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/plotcalc-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/style.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/intro/plotcalc.html
0.02Mb /work/scripting/doc/gnuplot/Kawano/datafile2-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/tics-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/misc2.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/index.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/label.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot3d.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/postscript-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot2-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/mo100.exp
0.05Mb /work/scripting/doc/gnuplot/Kawano/gallery/covar.dat
0.02Mb /work/scripting/doc/gnuplot/Kawano/gallery/covar.png
0.03Mb /work/scripting/doc/gnuplot/Kawano/gallery/wavefunc.dat
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/staircase.dat
0.24Mb /work/scripting/doc/gnuplot/Kawano/gallery/greenfunc.dat
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/nup.png
0.03Mb /work/scripting/doc/gnuplot/Kawano/gallery/integ2.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/overlap.dat
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/ddx15.dat
0.01Mb /work/scripting/doc/gnuplot/Kawano/gallery/twofig.dat
0.02Mb /work/scripting/doc/gnuplot/Kawano/gallery/twofig.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/fractal/selfsq1.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/fractal/selfsq2.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandelbrot0.png
0.05Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandelbrot1.png
0.04Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandelbrot2.png
0.03Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandelbrot3.png
0.08Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandelbrot4.png
0.03Mb /work/scripting/doc/gnuplot/Kawano/fractal/selfsquared1.png
0.07Mb /work/scripting/doc/gnuplot/Kawano/fractal/selfsquared2.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/fractal/mandel2.png
0.01Mb /work/scripting/doc/gnuplot/Kawano/index-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/set.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot6-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot1.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/datafile-e.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot2.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/tics.html
0.01Mb /work/scripting/doc/gnuplot/Kawano/plot6.html
0.38Mb /work/scripting/doc/gnuplot/gnuplot.html
0.82Mb /work/scripting/doc/gnuplot/gnuplot.ps
0.07Mb /work/scripting/doc/gnuplot/gnuplot-faq.html
0.05Mb /work/scripting/doc/python/fc/FPIG-paper.html
0.11Mb /work/scripting/doc/python/fc/pyfort_reference.htm
0.31Mb /work/scripting/doc/python/fc/pyfort_reference.pdf
0.03Mb /work/scripting/doc/python/fc/f2py-tutorial/eps/noise_zoom.eps
0.54Mb /work/scripting/doc/python/fc/f2py-tutorial/tutorial.pdf
0.01Mb /work/scripting/doc/python/fc/f2py-tutorial/tutorial_section1.tex
0.18Mb /work/scripting/doc/python/fc/f2py-tutorial/tutorial.ps.gz
0.01Mb /work/scripting/doc/python/fc/f2py-tutorial/lsodar/ClassIntegrate.py
0.09Mb /work/scripting/doc/python/fc/f2py-tutorial/lsodar/lsodar.f
0.10Mb /work/scripting/doc/python/fc/f2py.html
0.03Mb /work/scripting/doc/python/fc/swig_callback_ex/foo_wrap.c
0.01Mb /work/scripting/doc/python/PIL/decoder.html
0.02Mb /work/scripting/doc/python/PIL/image.html
0.02Mb /work/scripting/doc/python/PIL/intro01.html
0.01Mb /work/scripting/doc/python/PIL/formats.html
0.01Mb /work/scripting/doc/python/Pmw/PanedWidget.html
0.02Mb /work/scripting/doc/python/Pmw/MegaArchetype.html
0.02Mb /work/scripting/doc/python/Pmw/howtouse.html
0.01Mb /work/scripting/doc/python/Pmw/porting.html
0.01Mb /work/scripting/doc/python/Pmw/TimeCounter.html
0.01Mb /work/scripting/doc/python/Pmw/starting.html
0.01Mb /work/scripting/doc/python/Pmw/ButtonBox.html
0.01Mb /work/scripting/doc/python/Pmw/CounterDialog.html
0.01Mb /work/scripting/doc/python/Pmw/ComboBox.html
0.03Mb /work/scripting/doc/python/Pmw/PmwFunctions.html
0.01Mb /work/scripting/doc/python/Pmw/MessageBar.html
0.02Mb /work/scripting/doc/python/Pmw/HistoryText.html
0.02Mb /work/scripting/doc/python/Pmw/Counter.html
0.01Mb /work/scripting/doc/python/Pmw/bugs.html
0.01Mb /work/scripting/doc/python/Pmw/ScrolledText.html
0.01Mb /work/scripting/doc/python/Pmw/Color.html
0.01Mb /work/scripting/doc/python/Pmw/RadioSelect.html
0.04Mb /work/scripting/doc/python/Pmw/todo.html
0.01Mb /work/scripting/doc/python/Pmw/OptionMenu.html
0.01Mb /work/scripting/doc/python/Pmw/ScrolledCanvas.html
0.02Mb /work/scripting/doc/python/Pmw/MenuBar.html
0.02Mb /work/scripting/doc/python/Pmw/MainMenuBar.html
0.01Mb /work/scripting/doc/python/Pmw/MegaToplevel.html
0.02Mb /work/scripting/doc/python/Pmw/ScrolledFrame.html
0.02Mb /work/scripting/doc/python/Pmw/Balloon.html
0.01Mb /work/scripting/doc/python/Pmw/ScrolledText.gif
0.05Mb /work/scripting/doc/python/Pmw/changes.html
0.01Mb /work/scripting/doc/python/Pmw/NoteBook.html
0.02Mb /work/scripting/doc/python/Pmw/EntryField.html
0.01Mb /work/scripting/doc/python/Pmw/MessageDialog.html
0.01Mb /work/scripting/doc/python/Pmw/howtobuild.html
0.01Mb /work/scripting/doc/python/Pmw/ScrolledListBox.html
0.02Mb /work/scripting/doc/python/Tix/manpages/TixIntro.html
0.02Mb /work/scripting/doc/python/Tix/manpages/tixComboBox.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixScrolledListBox.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixTree.html
0.02Mb /work/scripting/doc/python/Tix/manpages/tixDisplayStyle.html
0.02Mb /work/scripting/doc/python/Tix/manpages/tixForm.html
0.02Mb /work/scripting/doc/python/Tix/manpages/tixGrid.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixFileEntry.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixExFileSelectBox.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixPanedWindow.html
0.06Mb /work/scripting/doc/python/Tix/manpages/tixHList.html
0.03Mb /work/scripting/doc/python/Tix/manpages/tixTList.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixListNoteBook.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixOptionMenu.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixSelect.html
0.01Mb /work/scripting/doc/python/Tix/manpages/compound.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixControl.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tix.html
0.01Mb /work/scripting/doc/python/Tix/manpages/tixNoteBook.html
0.08Mb /work/scripting/doc/python/Tix/pyguide.pdf
0.11Mb /work/scripting/doc/python/Tix/pytix.pdf
0.01Mb /work/scripting/doc/python/Tix/tix-book/fig/tlist/relation.gif
0.01Mb /work/scripting/doc/python/Tix/tix-book/fig/cover.gif
0.05Mb /work/scripting/doc/python/Tix/tix-book/fig/filesel/fb_comp.gif
0.02Mb /work/scripting/doc/python/Tix/tix-book/tlist.html
0.02Mb /work/scripting/doc/python/Tix/tix-book/container.html
0.03Mb /work/scripting/doc/python/Tix/tix-book/oop.html
0.01Mb /work/scripting/doc/python/Tix/tix-book/filesel.html
0.04Mb /work/scripting/doc/python/Tix/tix-book/intro.html
0.01Mb /work/scripting/doc/python/Tix/tix-book/hlist.html
0.04Mb /work/scripting/doc/python/unum/Unum_tutorial.html
0.04Mb /work/scripting/doc/python/jpython/review.html
0.01Mb /work/scripting/doc/python/jpython/faq.html
0.01Mb /work/scripting/doc/python/jpython/jpythonc.html
0.01Mb /work/scripting/doc/python/jpython/subclassing.html
0.02Mb /work/scripting/doc/python/jpython/JCPy-differences.html
0.01Mb /work/scripting/doc/python/jpython/usejava.html
0.03Mb /work/scripting/doc/python/spark.html
0.04Mb /work/scripting/doc/python/NumPy/Numeric/numpy.css
0.03Mb /work/scripting/doc/python/NumPy/Numeric/numpy-5.gif
0.04Mb /work/scripting/doc/python/NumPy/Numeric/numpy-12.html
0.03Mb /work/scripting/doc/python/NumPy/Numeric/numpy-13.html
0.04Mb /work/scripting/doc/python/NumPy/Numeric/numpy-14.html
0.01Mb /work/scripting/doc/python/NumPy/Numeric/numpy-17.html
0.01Mb /work/scripting/doc/python/NumPy/Numeric/numpy-18.html
0.02Mb /work/scripting/doc/python/NumPy/Numeric/numpy-19.html
0.12Mb /work/scripting/doc/python/NumPy/Numeric/numpy-22.html
0.01Mb /work/scripting/doc/python/NumPy/Numeric/numpy-5.html
0.07Mb /work/scripting/doc/python/NumPy/Numeric/numpy-6.html
0.03Mb /work/scripting/doc/python/NumPy/Numeric/numpy-7.html
0.05Mb /work/scripting/doc/python/NumPy/Numeric/numpy.html
0.05Mb /work/scripting/doc/python/NumPy/Numeric/numpy-9.html
0.05Mb /work/scripting/doc/python/NumPy/numeric_rewrite.pdf
1.23Mb /work/scripting/doc/python/NumPy/numpy.pdf
0.66Mb /work/scripting/doc/python/NumPy/NumTut/greece.pik
0.40Mb /work/scripting/doc/python/NumPy/numarray-0.5.pdf
0.40Mb /work/scripting/doc/python/NumPy/numarray-0.7.pdf
5.04Mb /work/scripting/doc/python/NumPy/numarray-0.5.ps
0.14Mb /work/scripting/doc/python/NumPy/numarray-0.7.html.tar.gz
0.01Mb /work/scripting/doc/python/NumPy/numarray/node53.html
0.05Mb /work/scripting/doc/python/NumPy/numarray/node58.html
0.03Mb /work/scripting/doc/python/NumPy/numarray/node60.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node61.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node6.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node65.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node21.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node22.html
0.03Mb /work/scripting/doc/python/NumPy/numarray/node23.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/contents.html
0.04Mb /work/scripting/doc/python/NumPy/numarray/genindex.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node30.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node31.html
0.04Mb /work/scripting/doc/python/NumPy/numarray/node33.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node34.html
0.01Mb /work/scripting/doc/python/NumPy/numarray/node37.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node38.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node39.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node41.html
0.02Mb /work/scripting/doc/python/NumPy/numarray/node42.html
0.28Mb /work/scripting/doc/python/NumPy/Asher_NumPy.html
0.04Mb /work/scripting/doc/python/SciPy/tutorial/img108.png
0.04Mb /work/scripting/doc/python/SciPy/tutorial/img109.png
0.01Mb /work/scripting/doc/python/SciPy/tutorial/images.tex
0.01Mb /work/scripting/doc/python/SciPy/tutorial/node8.html
0.03Mb /work/scripting/doc/python/SciPy/tutorial/images.pl
0.01Mb /work/scripting/doc/python/SciPy/tutorial/node21.html
0.01Mb /work/scripting/doc/python/SciPy/tutorial/node24.html
0.01Mb /work/scripting/doc/python/pymat/pymat.html
0.22Mb /work/scripting/doc/python/quickref2.1.html
0.06Mb /work/scripting/doc/python/quickref2.2/ar01s07.html
0.01Mb /work/scripting/doc/python/quickref2.2/ar01s08.html
0.01Mb /work/scripting/doc/python/quickref2.2/ar01s11.html
0.02Mb /work/scripting/doc/python/quickref2.2/ar01s12.html
0.02Mb /work/scripting/doc/python/quickref2.2/ar01s13.html
0.03Mb /work/scripting/doc/python/quickref2.2/ar01s16.html
0.01Mb /work/scripting/doc/python/quickref2.2/ar01s17.html
0.10Mb /work/scripting/doc/python/quickref2.2/ar01s18.html
0.24Mb /work/scripting/doc/python/quickref2.2/python22.pdf
0.01Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWeights.ps
0.02Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloBLT.ps
0.22Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWeights-pic.ps
0.02Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloMagnifier.ps
0.02Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWavesExt.ps
0.32Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloBLT-pic.ps
0.19Mb /work/scripting/doc/python/Pmw.Blt/ps/reference.ps
0.20Mb /work/scripting/doc/python/Pmw.Blt/ps/Pmw.Blt.doc.ps.gz
0.69Mb /work/scripting/doc/python/Pmw.Blt/ps/appetizer.ps
0.02Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWaves.ps
0.28Mb /work/scripting/doc/python/Pmw.Blt/ps/index.ps
0.03Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloUser.ps
1.01Mb /work/scripting/doc/python/Pmw.Blt/ps/tutorial.ps
0.01Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWorld2.ps
0.21Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloWorld1-pic.ps
0.45Mb /work/scripting/doc/python/Pmw.Blt/ps/HelloUser-pic.ps
0.10Mb /work/scripting/doc/python/Pmw.Blt/doc/reference.n
0.08Mb /work/scripting/doc/python/Pmw.Blt/doc/images/HelloWavesExt.gif
0.16Mb /work/scripting/doc/python/Pmw.Blt/doc/images/HelloVideo.gif
0.01Mb /work/scripting/doc/python/Pmw.Blt/doc/images/HelloMagnifier.gif
0.11Mb /work/scripting/doc/python/Pmw.Blt/doc/reference.html
0.02Mb /work/scripting/doc/python/Pmw.Blt/doc/tutorial.html
0.10Mb /work/scripting/doc/python/Pmw.Blt/doc/reference.sdf
0.01Mb /work/scripting/doc/python/Pmw.Blt/doc/python/html/HelloWavesExt.html
0.02Mb /work/scripting/doc/python/Pmw.Blt/doc/python/html/HelloUser.html
0.08Mb /work/scripting/doc/python/Pmw.Blt/private/reference.sdf.old
0.09Mb /work/scripting/doc/python/Pmw.Blt/private/input.sdf
0.01Mb /work/scripting/doc/python/Pmw.Blt/private/mail.0
0.01Mb /work/scripting/doc/python/Pmw.Blt/private/mail.2
0.15Mb /work/scripting/doc/python/Pmw.Blt/private/reference.html-orig
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/intObjects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/unicodeObjects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/sequence.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/fileObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/exceptions.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/mapping.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/profiling.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/importing.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/listObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/tupleObjects.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/arg-parsing.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/standardExceptions.html
0.06Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/type-structs.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/supporting-cycle-detection.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/bufferObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/unicodeMethodsAndSlots.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/stringObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/node81.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/node82.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/dictObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/refcountDetails.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/longObjects.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/object.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/exceptionHandling.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/builtinCodecs.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/threads.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/common-structs.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/allocating-objects.html
0.07Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/genindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/moduleObjects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/marshalling-utils.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/number.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/veryhigh.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/buffer-structs.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/api/initialization.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/info-units.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/inline-markup.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/directories.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/table-markup.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/latex-syntax.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/doc/indexing.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/errors.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/refcounts.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/node50.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/win-cookbook.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/callingPython.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/dnt-basics.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/using-cobjects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/node22.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/node23.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/node24.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ext/node32.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xml.sax.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-locale.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node374.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node689.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-pprint.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-weakref.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-posixfile.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xml.dom.minidom.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-fcntl.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/modindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/shlex-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-urlparse.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-audioop.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-string.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-signal.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-errno.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-email.Generator.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/obsolete-modules.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/condition-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/bltin-file-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node752.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/ossaudio-device-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node753.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-mailbox.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node126.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-email.Message.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-rfc822.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/audio-device-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node501.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/thread-objects.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/bytecodes.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-cd.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-cmath.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-socket.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/xdr-unpacker-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/other-gui-packages.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/form-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-codecs.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-htmllib.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-time.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/telnet-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-readline.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/python.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-process.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module--winreg.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/optparse-generating-help.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node509.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/nntp-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-asyncore.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-BaseHTTPServer.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-aifc.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node63.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node510.html
0.07Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/built-in-funcs.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-SocketServer.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-fd-ops.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/xmlparser-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-winsound.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-array.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/testresult-objects.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/curses-functions.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node268.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-webbrowser.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/match-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/SMTP-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node269.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/xdr-packer-objects.html
0.06Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/index.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-imageop.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xmlrpclib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/typesseq-mutable.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node270.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-file-dir.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/curses-textpad-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/zipfile-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node271.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/netdata.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/allos.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-random.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/formatter-interface.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-turtle.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-httplib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-types.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/set-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/ftp-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-pdb.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/typesseq-strings.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-thread.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xmllib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-math.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-sgmllib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node650.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/RawConfigParser-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/writer-interface.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node337.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-binascii.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-sys.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/string-methods.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/optparse-callback-examples.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-ConfigParser.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-email.Header.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/debugger-commands.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/pop3-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node281.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-chunk.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/message-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-urllib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node282.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/testcase-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xml.sax.handler.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/typesmapping.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-operator.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-newstreams.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/optparse-option-actions.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node658.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-threading.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node403.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/dom-node-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/imap4-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-curses.ascii.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-mpz.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node218.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-unicodedata.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/organizing-tests.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node406.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node720.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-HTMLParser.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-imp.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-path.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/tarfile-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-difflib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-traceback.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/MultiFile-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-fileinput.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/datetime-datetime.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/Cmd-objects.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/curses-window-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-imaplib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node293.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/datetime-time.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-textwrap.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-shutil.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-compiler.ast.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/datetime-tzinfo.html
0.05Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/contents.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/profile-stats.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-getopt.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-gc.html
0.06Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/lib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-tarfile.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/datetime-date.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/rexec-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-os.path.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/socket-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-stat.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node299.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/optparse-terminology.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/datetime-timedelta.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node545.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-logging.html
0.40Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/genindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-mimetypes.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/typesnumeric.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-zlib.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-nntplib.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/inspect-types.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-asynchat.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-bsddb.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-exceptions.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node105.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xml.sax.xmlreader.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-xml.dom.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-email.Charset.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-gl.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/content-handler-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/forms-objects.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/itertools-functions.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/typesseq.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-marshal.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/internet.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-stringprep.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/sequence-matcher.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/os-procinfo.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-struct.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/operator-map.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-email.Utils.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-mmap.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/node497.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/xmlreader-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-parser.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-rotor.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-calendar.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-tempfile.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/module-urllib2.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/dom-exceptions.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/re-syntax.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/lib/player-objects.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/modindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-macfs.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/mac.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-MacOS.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/toolbox.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/scripting.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/index.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-aepack.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-FrameWork.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/contents.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/node100.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/node101.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/genindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-aetypes.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/mac/module-EasyDialogs.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/numeric-types.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/function.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/naming.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/calls.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/try.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/index.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/assignment.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/import.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/slicings.html
0.05Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/types.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/contents.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/sequence-types.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/strings.html
0.08Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/genindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/node104.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/node105.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/comparisons.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/customization.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/ref.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/ref/binary.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node2.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node4.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node5.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node6.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node7.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node8.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node9.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/index.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node10.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node11.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node13.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node14.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/node15.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/tut/tut.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/module-distutils.sysconfig.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/postinstallation-script.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/simple-example.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/single-ext.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/source-dist.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/setup-config.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/dist/setup-script.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/inst/tweak-flags.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/inst/alt-install-windows.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/inst/config-syntax.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/inst/standard-install.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/inst/search-path.html
0.03Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/modindex.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/whatsnew/section-generators.html
0.02Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/whatsnew/node17.html
0.04Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/whatsnew/node18.html
0.01Mb /work/scripting/doc/python/Reference/Python-Docs-2.3/whatsnew/node20.html
0.01Mb /work/scripting/doc/python/parallel/pypar.txt
0.07Mb /work/scripting/doc/python/parallel/parallel_python.pdf
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/NavigableTree_NavigableTree.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/Table_Column.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/ConnectedBox_ConnectedBox.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/ShadowBox_ShadowBox.py.html
0.04Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/GuiAppD_GuiAppD.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Client/wcc_protocol_WackyConnection.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Client/wcc_dialog_MessageDialog.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Client/wcc_client_Hermes.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Server/wimd_pwfile_wimd_pwfile.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Server/wimd_server_wimd_channel.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Server/wimd_server_wimd_server.py.html
0.03Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/SampleApps/WhackyChat/Server/CommandLineApp_CommandLineApp.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/AnimatedFileIcon_AnimatedFileIcon.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/PipeOutputWindow_PipeOutputWindow.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/AnimatedFolder_FileFolder.py.html
0.03Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/UserPrefs_UserPrefs.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/ProgressMeter_ProgressMeter.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/AnimatedIcon_AnimatedIcon.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/TreeNavigator_TreeNavigator.py.html
0.01Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/FontChooserDialog_FontChooserDialog.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/PmwContribD-r2_0_1/StructuredText.py.html
0.02Mb /work/scripting/doc/python/PmwContribD/index.html
0.01Mb /work/scripting/doc/python/dislin/disipyl/tutorial.html
0.02Mb /work/scripting/doc/python/happydoc/doc/index.html
0.02Mb /work/scripting/doc/python/happydoc/README.txt
0.21Mb /work/scripting/doc/python/py-in-10pages.ps
0.01Mb /work/scripting/doc/python/pybliographer/documentation/main.png
0.14Mb /work/scripting/doc/python/quickref2.1.txt
0.24Mb /work/scripting/doc/python/quickref2.2.pdf
0.02Mb /work/scripting/doc/python/Py_vs_Perl_vs_Tcl.txt
0.02Mb /work/scripting/doc/python/Scientific-Python/html/Scientific_25.html
0.01Mb /work/scripting/doc/python/Scientific-Python/html/Scientific_3.html
0.32Mb /work/scripting/doc/python/Scientific-Python/manual.pdf
0.10Mb /work/scripting/doc/python/Scientific-Python/SciComp-wPython.ps
0.01Mb /work/scripting/doc/python/Tkinter/life-preserver/ClassText.html
0.01Mb /work/scripting/doc/python/Tkinter/life-preserver/ClassCanvas.html
0.02Mb /work/scripting/doc/python/Tkinter/intro/dialog-windows.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/x1366-options.htm
0.02Mb /work/scripting/doc/python/Tkinter/intro/canvasarc1.gif
0.02Mb /work/scripting/doc/python/Tkinter/intro/x1728-methods.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/x6637-options.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/x9170-window-related-information.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/x8518-options.htm
0.03Mb /work/scripting/doc/python/Tkinter/intro/WindowsFonts.gif
0.03Mb /work/scripting/doc/python/Tkinter/intro/x7991-methods.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/SystemFonts.gif
0.02Mb /work/scripting/doc/python/Tkinter/intro/BuiltinCursors.gif
0.01Mb /work/scripting/doc/python/Tkinter/intro/grid3.gif
0.01Mb /work/scripting/doc/python/Tkinter/intro/index.htm
0.02Mb /work/scripting/doc/python/Tkinter/intro/x7505-concepts.htm
0.01Mb /work/scripting/doc/python/Tkinter/intro/x3565-options.htm
0.02Mb /work/scripting/doc/python/Tkinter/intro/events-and-bindings.htm
0.02Mb /work/scripting/doc/python/Tkinter/intro/canvasbitmap1.gif
0.01Mb /work/scripting/doc/python/Tkinter/intro/x444-fonts.htm
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassText.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassCanvas.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassMenubutton.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassRadiobutton.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassToplevel.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassMenu.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassCheckbutton.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassButton.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassScale.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassListbox.html
0.01Mb /work/scripting/doc/python/Tkinter/manpages/ClassEntry.html
0.39Mb /work/scripting/doc/python/Tkinter/quickref-Tkinter.pdf
0.13Mb /work/scripting/doc/python/biggles/libplot_C.html
0.01Mb /work/scripting/doc/python/biggles/refmanual/components.html
0.01Mb /work/scripting/doc/python/optimize-python.html
0.02Mb /work/scripting/doc/python/styleguide/docstring-style.html
0.03Mb /work/scripting/doc/python/styleguide/Py-style.html
0.01Mb /work/scripting/doc/python/Gnuplot/doc/index.html
0.03Mb /work/scripting/doc/python/Gnuplot/doc/_Gnuplot.py_Gnuplot.html
0.01Mb /work/scripting/doc/python/Gnuplot/doc/PlotItems.py_PlotItem.html
0.03Mb /work/scripting/doc/python/Gnuplot/doc/Gnuplot/_Gnuplot.py_Gnuplot.html
0.01Mb /work/scripting/doc/python/Gnuplot/doc/Gnuplot/PlotItems.py_PlotItem.html
0.01Mb /work/scripting/doc/python/Gnuplot/index.html
0.03Mb /work/scripting/doc/python/Gnuplot/_Gnuplot.py_Gnuplot.html
0.01Mb /work/scripting/doc/python/Gnuplot/PlotItems.py_PlotItem.html
0.03Mb /work/scripting/doc/python/Gnuplot/Gnuplot/_Gnuplot.py_Gnuplot.html
0.01Mb /work/scripting/doc/python/Gnuplot/Gnuplot/PlotItems.py_PlotItem.html
0.37Mb /work/scripting/doc/python/Python-FAQ.html
0.05Mb /work/scripting/doc/python/IDLE-doc/idle2.html
/work/scripting/doc/python/NumPy/numarray-0.5.ps 5.04Mb
/work/scripting/doc/latex/intro/teTeX/latex/graphics/epslatex.ps 2.31Mb
/work/scripting/doc/latex/intro/teTeX/generic/xypic/xyrefer.ps 1.86Mb
/work/scripting/doc/python/Pmw.Blt/ps/tutorial.ps 1.01Mb


version 3 of tree traversal: root= /work/scripting/doc
1.01Mb file in /work/scripting/doc/latex/intro/ltxprimer-1.0.pdf
1.31Mb file in /work/scripting/doc/latex/intro/tipaman.pdf
0.77Mb file in /work/scripting/doc/latex/intro/epslatex.ps
1.39Mb file in /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctfull.html
2.82Mb file in /work/scripting/doc/latex/intro/teTeX/context/base/ms-cb-en.pdf
0.79Mb file in /work/scripting/doc/latex/intro/teTeX/metapost/base/mpman.ps
2.31Mb file in /work/scripting/doc/latex/intro/teTeX/latex/graphics/epslatex.ps
0.98Mb file in /work/scripting/doc/latex/intro/teTeX/generic/pstricks/doc-fill.ps
0.67Mb file in /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyguide.ps
1.86Mb file in /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyrefer.ps
0.82Mb file in /work/scripting/doc/gnuplot/gnuplot.ps
0.54Mb file in /work/scripting/doc/python/fc/f2py-tutorial/tutorial.pdf
1.23Mb file in /work/scripting/doc/python/NumPy/numpy.pdf
5.04Mb file in /work/scripting/doc/python/NumPy/numarray-0.5.ps
0.66Mb file in /work/scripting/doc/python/NumPy/NumTut/greece.pik
0.69Mb file in /work/scripting/doc/python/Pmw.Blt/ps/appetizer.ps
1.01Mb file in /work/scripting/doc/python/Pmw.Blt/ps/tutorial.ps
creating mynewdir
removing mynewdir
You have a non-existing directory
    /work/maple/bin 
in your path
You have a non-existing directory
    /work/matlab/bin 
in your path
You have a non-existing directory
    /local/TEX/bin.linux 
in your path
You have a non-existing directory
    /work/maple7/bin 
in your path
You have a non-existing directory
    /work/NO/la/bin/Linux/opt 
in your path
You have a non-existing directory
    /work/sysdir/src/java/jdk1.3/bin 
in your path
You have a non-existing directory
    /usr/local/FFC/bin 
in your path
vtk  not found
leading text ['listitem1', 'listitem2']
another leading text ['listitem1', 'listitem2']
No leading text ['listitem1', 'listitem2']
No leading text /home/hpl
statistics: avg=$avg, min=$min, max=$max

before swap: v1= 1.3  v2= some text
after  swap: v1= 1.3  v2= some text
files of *.ps *.gif and *.py type:
tmp_c_runs.ps
tmp.ps
tmp_c.gif
NumPy_basics.py
hw.py
leastsquares.py
Grid2D.py
datatrans1.py
datatrans2.py
ScientificPython.py
datatrans-eff.py
datatrans3a.py
datatrans3b.py
datatrans3c.py
datatrans3d.py
loop4simviz1.py
loop4simviz2.py
tmp.py
commontasks.py
simviz1.py
simviz2.py
convert1.py
convert2.py
SciPy.py
Output of the command perl -pe '' hw.py was

#!/usr/bin/env python
import sys, math       # load system and math module
r = float(sys.argv[1]) # extract the 1st command-line arg.
s = math.sin(r)
print "Hello, World! sin(" + str(r) + ")=" + str(s)
file= /usr/home/hpl/scripting/perl/intro/hw.pl
head= /usr/home/hpl/scripting/perl/intro
tail= hw.pl
dirname = /usr/home/hpl/scripting/perl/intro
basename= hw.pl

Yes! created tmp/some/tmp/tmp


Programming with classes:
MyBase: i= 5 j= 7
MySub: i= 7 j= 8 k= 9
i1 is MyBase
i2 is MySub
i2 is MyBase too
i1.__dict__: {'i': 5, 'j': 7}
i2.__dict__: {'i': 7, 'k': 9, 'j': 8}
Names: MyBase MyBase.write
dir(i1): ['__doc__', '__init__', '__module__', 'i', 'j', 'write']
dir(i2): ['__doc__', '__init__', '__module__', 'i', 'j', 'k', 'write']
some string
['__doc__', '__init__', '__module__', 'i', 'j', 'k', 'q', 'write']



list[6] raises an exception
Exception type= exceptions.IndexError
Exception value= list index out of range
average= 2.0
average= Empty argument list in average
Exception type= Empty argument list in average
Exception value= None
Exception type= exceptions.IOError
Exception value= [Errno 2] No such file or directory: 'ppp'
item 0: -                     description: initial shape of u
item 1: t                     description: initial shape of H
item 2: s                     description: shape of u at time=2.5
curve1                description: initial shape of u
curve2                description: initial shape of H
curve3                description: shape of u at time=2.5
1.2 is greater than or equal to 100 (a is <type 'str'> and b is <type 'int'> )
1.2 is less than 100 (a is <type 'float'> and b is <type 'int'> )
testing string b < 100: error!
testing float(b) < 100: ok
{
   'A' : [1.2, -3.3999999999999999, 5.5, -9, 100],
   'INDENT' : 2,
   'MyBase' : <class __main__.MyBase at 0x4081889c>,
   'MySub' : <class __main__.MySub at 0x408188cc>,
   '__builtins__' : <module '__builtin__' (built-in)>,
   '__doc__' : ':"\nexec python $0 ${1+"$@"}\n',
   '__file__' : './commontasks.py',
   '__name__' : '__main__',
   '__warningregistry__' : {
       ('raising a string exception is deprecated', <class exceptions.PendingDeprecationWarning at 0x401dbf2c>, 444) : 1,
       },
   'a' : 0.59999999999999998,
   'api_version' : 1012,
   'arg_counter' : 6,
   'arglist' : ['myarg1', 'displacement', 'tmp.ps', 'myvar2'],
   'argv' : ['./commontasks.py'],
   'average' : <function average at 0x40823a74>,
   'average_exc' : 'Empty argument list in average',
   'avg' : 4.2249999999999996,
   'b' : '1.2',
   'basename' : 'hw.pl',
   'bigfiles' : ['1.01Mb file in /work/scripting/doc/latex/intro/ltxprimer-1.0.pdf', '1.31Mb file in /work/scripting/doc/latex/intro/tipaman.pdf', '0.77Mb file in /work/scripting/doc/latex/intro/epslatex.ps', '1.39Mb file in /work/scripting/doc/latex/intro/teTeX/help/Catalogue/ctfull.html', '2.82Mb file in /work/scripting/doc/latex/intro/teTeX/context/base/ms-cb-en.pdf', '0.79Mb file in /work/scripting/doc/latex/intro/teTeX/metapost/base/mpman.ps', '2.31Mb file in /work/scripting/doc/latex/intro/teTeX/latex/graphics/epslatex.ps', '0.98Mb file in /work/scripting/doc/latex/intro/teTeX/generic/pstricks/doc-fill.ps', '0.67Mb file in /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyguide.ps', '1.86Mb file in /work/scripting/doc/latex/intro/teTeX/generic/xypic/xyrefer.ps', '0.82Mb file in /work/scripting/doc/gnuplot/gnuplot.ps', '0.54Mb file in /work/scripting/doc/python/fc/f2py-tutorial/tutorial.pdf', '1.23Mb file in /work/scripting/doc/python/NumPy/numpy.pdf', '5.04Mb file in /work/scripting/doc/python/NumPy/numarray-0.5.ps', '0.66Mb file in /work/scripting/doc/python/NumPy/NumTut/greece.pik', '0.69Mb file in /work/scripting/doc/python/Pmw.Blt/ps/appetizer.ps', '1.01Mb file in /work/scripting/doc/python/Pmw.Blt/ps/tutorial.ps'],
   'builtin_module_names' : ('__builtin__', '__main__', '_codecs', '_sre', '_symtable', 'errno', 'exceptions', 'gc', 'imp', 'marshal', 'posix', 'signal', 'sys', 'thread', 'xxsubtype', 'zipimport'),
   'byteorder' : 'little',
   'call_tracing' : <built-in function call_tracing>,
   'callstats' : <built-in function callstats>,
   'checksize1' : <function checksize1 at 0x408235a4>,
   'checksize2' : <function checksize2 at 0x4023772c>,
   'checksize3' : <function checksize3 at 0x40823064>,
   'cmd' : "perl -pe '' hw.py",
   'cmlargs' : {
       '-c_in_H' : '9.8',
       '-tstop' : '6.1',
       },
   'compare' : <function compare at 0x40823b54>,
   'copyright' : 'Copyright (c) 2001, 2002, 2003 Python Software Foundation.\nAll Rights Reserved.\n\nCopyright (c) 2000 BeOpen.com.\nAll Rights Reserved.\n\nCopyright (c) 1995-2001 Corporation for National Research Initiatives.\nAll Rights Reserved.\n\nCopyright (c) 1991-1995 Stichting Mathematisch Centrum, Amsterdam.\nAll Rights Reserved.',
   'curvelist' : [('curve1', 'initial shape of u'), ('curve2', 'initial shape of H'), ('curve3', 'shape of u at time=2.5')],
   'd' : '.',
   'directory' : 'tmp/some/tmp/tmp',
   'dirname' : '/usr/home/hpl/scripting/perl/intro',
   'displayhook' : <built-in function displayhook>,
   'displaylist' : <function displaylist at 0x40823ae4>,
   'displaylist2' : <function displaylist2 at 0x40823b1c>,
   'dump1' : <function dump1 at 0x40823614>,
   'dump2' : <function dump2 at 0x4082364c>,
   'entry' : 1073569782,
   'exc_clear' : <built-in function exc_clear>,
   'exc_info' : <built-in function exc_info>,
   'exc_traceback' : <traceback object at 0x408217fc>,
   'exc_type' : <class exceptions.IOError at 0x401db47c>,
   'exc_value' : <exceptions.IOError instance at 0x408282ac>,
   'excepthook' : <built-in function excepthook>,
   'exec_prefix' : '/usr',
   'executable' : '/usr/bin/python',
   'exit' : <built-in function exit>,
   'exitfunc' : <function _run_exitfuncs at 0x4024f6bc>,
   'explanations' : ['initial shape of u', 'initial shape of H', 'shape of u at time=2.5'],
   'file' : 'SciPy.py',
   'fileinfo' : '1.01Mb file in /work/scripting/doc/python/Pmw.Blt/ps/tutorial.ps',
   'filelist' : ['NumPy_basics.py', 'hw.py', 'leastsquares.py', 'Grid2D.py', 'datatrans1.py', 'datatrans2.py', 'ScientificPython.py', 'datatrans-eff.py', 'datatrans3a.py', 'datatrans3b.py', 'datatrans3c.py', 'datatrans3d.py', 'loop4simviz1.py', 'loop4simviz2.py', 'tmp.py', 'commontasks.py', 'simviz1.py', 'simviz2.py', 'convert1.py', 'convert2.py', 'SciPy.py'],
   'filename' : 'hw.py',
   'filesize' : 202L,
   'filesort' : <function filesort at 0x4082341c>,
   'find' : <function find at 0x4081ebfc>,
   'fnmatch' : <module 'fnmatch' from '/usr/lib/python2.3/fnmatch.pyc'>,
   'found' : 0,
   'getcheckinterval' : <built-in function getcheckinterval>,
   'getdefaultencoding' : <built-in function getdefaultencoding>,
   'getdlopenflags' : <built-in function getdlopenflags>,
   'getfilesystemencoding' : <built-in function getfilesystemencoding>,
   'getrecursionlimit' : <built-in function getrecursionlimit>,
   'getrefcount' : <built-in function getrefcount>,
   'glob' : <module 'glob' from '/usr/lib/python2.3/glob.pyc'>,
   'head' : '/usr/home/hpl/scripting/perl/intro',
   'here' : '/home/work/scripting/src/py/intro',
   'hexversion' : 33752048,
   'i' : 4,
   'i1' : <__main__.MyBase instance at 0x4081bf2c>,
   'i2' : <__main__.MySub instance at 0x4081ba6c>,
   'infile' : <closed file '.myprog.cpp', mode 'r' at 0x4045cae0>,
   'infilename' : '.myprog.cpp',
   'item' : '-tstop',
   'last_access' : 1079261774,
   'line' : 'print "Hello, World! sin(" + str(r) + ")=" + str(s)\n',
   'line1' : 'iteration 12:    eps= 1.245E-05',
   'line2' : '.myc_12@displacement@u(x,3.1415)@  no upwinding',
   'line_no' : 7,
   'lines' : ['#!/usr/bin/env python\n', 'import sys, math       # load system and math module\n', 'r = float(sys.argv[1]) # extract the 1st command-line arg.\n', 's = math.sin(r)\n', 'print "Hello, World! sin(" + str(r) + ")=" + str(s)\n'],
   'list' : ['t1', 't2', 't3'],
   'math' : <module 'math' from '/usr/lib/python2.3/lib-dynload/math.so'>,
   'max' : 9,
   'maxint' : 2147483647,
   'maxunicode' : 1114111,
   'meta_path' : [],
   'min' : 1,
   'mode' : 33261,
   'modules' : {
       'ArrayPrinter' : <module 'ArrayPrinter' from '/usr/lib/python2.3/site-packages/Numeric/ArrayPrinter.pyc'>,
       'Gnuplot' : <module 'Gnuplot' from '/home/hpl/install/lib/python/Gnuplot/__init__.pyc'>,
       'Gnuplot.Numeric' : None,
       'Gnuplot.PlotItems' : <module 'Gnuplot.PlotItems' from '/home/hpl/install/lib/python/Gnuplot/PlotItems.pyc'>,
       'Gnuplot._Gnuplot' : <module 'Gnuplot._Gnuplot' from '/home/hpl/install/lib/python/Gnuplot/_Gnuplot.pyc'>,
       'Gnuplot.cStringIO' : None,
       'Gnuplot.gp' : <module 'Gnuplot.gp' from '/home/hpl/install/lib/python/Gnuplot/gp.pyc'>,
       'Gnuplot.gp_unix' : <module 'Gnuplot.gp_unix' from '/home/hpl/install/lib/python/Gnuplot/gp_unix.pyc'>,
       'Gnuplot.os' : None,
       'Gnuplot.string' : None,
       'Gnuplot.sys' : None,
       'Gnuplot.tempfile' : None,
       'Gnuplot.utils' : <module 'Gnuplot.utils' from '/home/hpl/install/lib/python/Gnuplot/utils.pyc'>,
       'Numeric' : <module 'Numeric' from '/usr/lib/python2.3/site-packages/Numeric/Numeric.pyc'>,
       'Pmw' : <Pmw.Pmw_1_2.lib.PmwLoader.PmwLoader instance at 0x402557cc>,
       'Pmw.Pmw_1_2' : <module 'Pmw.Pmw_1_2' from '/work/sysdir/src/python/tools/Pmw/Pmw_1_2/__init__.pyc'>,
       'Pmw.Pmw_1_2.lib' : <module 'Pmw.Pmw_1_2.lib' from '/work/sysdir/src/python/tools/Pmw/Pmw_1_2/lib/__init__.pyc'>,
       'Pmw.Pmw_1_2.lib.PmwLoader' : <module 'Pmw.Pmw_1_2.lib.PmwLoader' from '/work/sysdir/src/python/tools/Pmw/Pmw_1_2/lib/PmwLoader.pyc'>,
       'Pmw.Pmw_1_2.lib.os' : None,
       'Pmw.Pmw_1_2.lib.string' : None,
       'Pmw.Pmw_1_2.lib.sys' : None,
       'Pmw.Pmw_1_2.lib.types' : None,
       'Pmw.os' : None,
       'Pmw.re' : None,
       'Pmw.sys' : None,
       'Precision' : <module 'Precision' from '/usr/lib/python2.3/site-packages/Numeric/Precision.pyc'>,
       'StringIO' : <module 'StringIO' from '/usr/lib/python2.3/StringIO.pyc'>,
       'Tkconstants' : <module 'Tkconstants' from '/usr/lib/python2.3/lib-tk/Tkconstants.pyc'>,
       'Tkinter' : <module 'Tkinter' from '/usr/lib/python2.3/lib-tk/Tkinter.pyc'>,
       'UserDict' : <module 'UserDict' from '/usr/lib/python2.3/UserDict.pyc'>,
       '_Pmw' : <module 'Pmw' from '/work/sysdir/src/python/tools/Pmw/__init__.pyc'>,
       '__builtin__' : <module '__builtin__' (built-in)>,
       '__future__' : <module '__future__' from '/usr/lib/python2.3/__future__.pyc'>,
       '__main__' : <module '__main__' from './commontasks.py'>,
       '_codecs' : <module '_codecs' (built-in)>,
       '_dotblas' : <module '_dotblas' from '/usr/lib/python2.3/site-packages/Numeric/_dotblas.so'>,
       '_iconv_codec' : <module '_iconv_codec' from '/usr/lib/python2.3/site-packages/_iconv_codec.so'>,
       '_numpy' : <module '_numpy' from '/usr/lib/python2.3/site-packages/Numeric/_numpy.so'>,
       '_random' : <module '_random' from '/usr/lib/python2.3/lib-dynload/_random.so'>,
       '_sre' : <module '_sre' (built-in)>,
       '_tkinter' : <module '_tkinter' from '/usr/lib/python2.3/lib-dynload/_tkinter.so'>,
       'atexit' : <module 'atexit' from '/usr/lib/python2.3/atexit.pyc'>,
       'binascii' : <module 'binascii' from '/usr/lib/python2.3/lib-dynload/binascii.so'>,
       'cStringIO' : <module 'cStringIO' from '/usr/lib/python2.3/lib-dynload/cStringIO.so'>,
       'codecs' : <module 'codecs' from '/usr/lib/python2.3/codecs.pyc'>,
       'copy' : <module 'copy' from '/usr/lib/python2.3/copy.pyc'>,
       'copy_reg' : <module 'copy_reg' from '/usr/lib/python2.3/copy_reg.pyc'>,
       'dotblas' : <module 'dotblas' from '/usr/lib/python2.3/site-packages/Numeric/dotblas/__init__.pyc'>,
       'dotblas.Numeric' : None,
       'dotblas._dotblas' : None,
       'dotblas._numpy' : None,
       'dotblas.multiarray' : None,
       'encodings' : <module 'encodings' from '/usr/lib/python2.3/encodings/__init__.pyc'>,
       'encodings.aliases' : <module 'encodings.aliases' from '/usr/lib/python2.3/encodings/aliases.pyc'>,
       'encodings.codecs' : None,
       'encodings.encodings' : None,
       'encodings.exceptions' : None,
       'encodings.latin_1' : <module 'encodings.latin_1' from '/usr/lib/python2.3/encodings/latin_1.pyc'>,
       'encodings.types' : None,
       'errno' : <module 'errno' (built-in)>,
       'exceptions' : <module 'exceptions' (built-in)>,
       'fcntl' : <module 'fcntl' from '/usr/lib/python2.3/lib-dynload/fcntl.so'>,
       'fnmatch' : <module 'fnmatch' from '/usr/lib/python2.3/fnmatch.pyc'>,
       'getopt' : <module 'getopt' from '/usr/lib/python2.3/getopt.pyc'>,
       'glob' : <module 'glob' from '/usr/lib/python2.3/glob.pyc'>,
       'iconv_codec' : <module 'iconv_codec' from '/usr/lib/python2.3/site-packages/iconv_codec.pyc'>,
       'linecache' : <module 'linecache' from '/usr/lib/python2.3/linecache.pyc'>,
       'marshal' : <module 'marshal' (built-in)>,
       'math' : <module 'math' from '/usr/lib/python2.3/lib-dynload/math.so'>,
       'multiarray' : <module 'multiarray' from '/usr/lib/python2.3/site-packages/Numeric/multiarray.so'>,
       'numeric_version' : <module 'numeric_version' from '/usr/lib/python2.3/site-packages/Numeric/numeric_version.pyc'>,
       'os' : <module 'os' from '/usr/lib/python2.3/os.pyc'>,
       'os.path' : <module 'posixpath' from '/usr/lib/python2.3/posixpath.pyc'>,
       'pickle' : <module 'pickle' from '/usr/lib/python2.3/pickle.pyc'>,
       'posix' : <module 'posix' (built-in)>,
       'posixpath' : <module 'posixpath' from '/usr/lib/python2.3/posixpath.pyc'>,
       'py4cs' : <module 'py4cs' from '/work/scripting/src/tools/py4cs/__init__.pyc'>,
       'py4cs.FuncDependenceViz' : <module 'py4cs.FuncDependenceViz' from '/work/scripting/src/tools/py4cs/FuncDependenceViz.pyc'>,
       'py4cs.Gnuplot' : None,
       'py4cs.Numeric' : None,
       'py4cs.Pmw' : None,
       'py4cs.Tkinter' : None,
       'py4cs.funcs' : <module 'py4cs.funcs' from '/work/scripting/src/tools/py4cs/funcs.pyc'>,
       'py4cs.getopt' : None,
       'py4cs.math' : None,
       'py4cs.os' : None,
       'py4cs.re' : None,
       'py4cs.shutil' : None,
       'py4cs.sys' : None,
       'py4cs.threading' : None,
       'py4cs.time' : None,
       'random' : <module 'random' from '/usr/lib/python2.3/random.pyc'>,
       're' : <module 're' from '/usr/lib/python2.3/re.pyc'>,
       'shutil' : <module 'shutil' from '/usr/lib/python2.3/shutil.pyc'>,
       'signal' : <module 'signal' (built-in)>,
       'site' : <module 'site' from '/usr/lib/python2.3/site.pyc'>,
       'sre' : <module 'sre' from '/usr/lib/python2.3/sre.pyc'>,
       'sre_compile' : <module 'sre_compile' from '/usr/lib/python2.3/sre_compile.pyc'>,
       'sre_constants' : <module 'sre_constants' from '/usr/lib/python2.3/sre_constants.pyc'>,
       'sre_parse' : <module 'sre_parse' from '/usr/lib/python2.3/sre_parse.pyc'>,
       'stat' : <module 'stat' from '/usr/lib/python2.3/stat.pyc'>,
       'string' : <module 'string' from '/usr/lib/python2.3/string.pyc'>,
       'strop' : <module 'strop' from '/usr/lib/python2.3/lib-dynload/strop.so'>,
       'struct' : <module 'struct' from '/usr/lib/python2.3/lib-dynload/struct.so'>,
       'sys' : <module 'sys' (built-in)>,
       'tempfile' : <module 'tempfile' from '/usr/lib/python2.3/tempfile.pyc'>,
       'thread' : <module 'thread' (built-in)>,
       'threading' : <module 'threading' from '/usr/lib/python2.3/threading.pyc'>,
       'time' : <module 'time' from '/usr/lib/python2.3/lib-dynload/time.so'>,
       'traceback' : <module 'traceback' from '/usr/lib/python2.3/traceback.pyc'>,
       'types' : <module 'types' from '/usr/lib/python2.3/types.pyc'>,
       'umath' : <module 'umath' from '/usr/lib/python2.3/site-packages/Numeric/umath.so'>,
       'warnings' : <module 'warnings' from '/usr/lib/python2.3/warnings.pyc'>,
       'zipimport' : <module 'zipimport' (built-in)>,
       },
   'myarg1' : 'myarg1',
   'myargs' : ['-myopt', '9.9', '-tstop', '6.1', '-c_in_H', '9.8'],
   'myfile' : 'hw.py',
   'myfile_stat' : (33261, 68938L, 778L, 1, 8029, 8029, 202L, 1079261774, 1071617117, 1073569782),
   'myvar2' : 'myvar2',
   'name' : '/usr/home/hpl/scripting/perl/intro/hw.pl',
   'newline1' : 'iteration#12:#eps=#1.245E-05',
   'option' : '-c_in_H',
   'os' : <module 'os' from '/usr/lib/python2.3/os.pyc'>,
   'outfile' : <open file '.myprog2.cpp', mode 'a' at 0x40230c20>,
   'outfilename' : '.myprog2.cpp',
   'path' : ['/home/work/scripting/src/py/intro', '/home/hpl/hp/div/Ola-install', '/work/sysdir/Linux/lib/vtk', '/work/sysdir/src/VTK/Wrapping/Python', '/work/sysdir/Linux/dislin/python', '/home/hpl/install/lib/python', '/work/sysdir/src/python/tools', '/work/sysdir/src/python/lib', '/work/scripting/src/tools', '/work/sysdir/src/python/Python-2.3/Tools', '/home/work/scripting/src/py/intro', '/home/hpl/hp/pyPDE/src/lib', '/home/hpl/hp/pyPDE/src/lib/idlelib', '/work/NO/bin', '/usr/lib/python23.zip', '/usr/lib/python2.3', '/usr/lib/python2.3/plat-linux2', '/usr/lib/python2.3/lib-tk', '/usr/lib/python2.3/lib-dynload', '/usr/local/lib/python2.3/site-packages', '/usr/lib/python2.3/site-packages', '/usr/lib/python2.3/site-packages/HTMLgen', '/usr/lib/python2.3/site-packages/Numeric', '/usr/lib/python2.3/site-packages/PIL', '/usr/lib/python2.3/site-packages/gtk-2.0', '/usr/lib/python2.3/site-packages/vtk_python', '/usr/lib/site-python'],
   'path_hooks' : [<type 'zipimport.zipimporter'>],
   'path_importer_cache' : {
       '' : None,
       '/home/hpl/hp/div/Ola-install' : None,
       '/home/hpl/hp/pyPDE/src/lib' : None,
       '/home/hpl/hp/pyPDE/src/lib/idlelib' : None,
       '/home/hpl/install/lib/python' : None,
       '/home/hpl/install/lib/python/Gnuplot' : None,
       '/home/work/scripting/src/py/intro' : None,
       '/usr/lib/python2.3' : None,
       '/usr/lib/python2.3/' : None,
       '/usr/lib/python2.3/encodings' : None,
       '/usr/lib/python2.3/lib-dynload' : None,
       '/usr/lib/python2.3/lib-tk' : None,
       '/usr/lib/python2.3/plat-linux2' : None,
       '/usr/lib/python2.3/site-packages' : None,
       '/usr/lib/python2.3/site-packages/HTMLgen' : None,
       '/usr/lib/python2.3/site-packages/Numeric' : None,
       '/usr/lib/python2.3/site-packages/Numeric/dotblas' : None,
       '/usr/lib/python2.3/site-packages/PIL' : None,
       '/usr/lib/python2.3/site-packages/gtk-2.0' : None,
       '/usr/lib/python2.3/site-packages/vtk_python' : None,
       '/usr/lib/python23.zip' : None,
       '/usr/lib/site-python' : None,
       '/usr/local/lib/python2.3/site-packages' : None,
       '/work/NO/bin' : None,
       '/work/scripting/src/tools' : None,
       '/work/scripting/src/tools/py4cs' : None,
       '/work/sysdir/Linux/dislin/python' : None,
       '/work/sysdir/Linux/lib/vtk' : None,
       '/work/sysdir/src/VTK/Wrapping/Python' : None,
       '/work/sysdir/src/python/Python-2.3/Tools' : None,
       '/work/sysdir/src/python/lib' : None,
       '/work/sysdir/src/python/tools' : None,
       '/work/sysdir/src/python/tools/Pmw' : None,
       '/work/sysdir/src/python/tools/Pmw/Pmw_1_2' : None,
       '/work/sysdir/src/python/tools/Pmw/Pmw_1_2/lib' : None,
       },
   'paths' : ['/home/hpl/bin', '/work/maple/bin', '/work/matlab/bin', '/local/TEX/bin.linux', '/work/scripting/src/tools', '/work/scripting/Linux/bin', '/bin', '/usr/bin', '/usr/X11R6/bin', '/usr/sbin', '/work/maple7/bin', '/home/hpl/install/bin', '/home/hpl/hp/pyPDE/src/lib', '/work/NO/bin', '/work/NO/md/bin/Linux/opt', '/work/NO/dp/bin/Linux/opt', '/work/NO/bt/bin/Linux/opt', '/work/NO/la/bin/Linux/opt', '/work/sysdir/Linux/bin', '/work/NO/internal/bin', '/usr/local/Acrobat5/bin', '/work/sysdir/src/java/jdk1.3/bin', '/work/sysdir/src/python/Jython/jython-2.0', '/usr/local/FFC/bin', '.'],
   'pipe' : <closed file 'sh', mode 'w' at 0x402302a0>,
   'platform' : 'linux2',
   'plottitle' : 'displacement',
   'prefix' : '/usr',
   'pretty_dict_print' : <function pretty_dict_print at 0x40823b8c>,
   'program' : 'vtk',
   'psfile' : 'tmp.ps',
   'r' : 100,
   're' : <module 're' from '/usr/lib/python2.3/re.pyc'>,
   'regex' : <_sre.SRE_Match object at 0x4022eaa0>,
   'res' : ['#!/usr/bin/env python\n', 'import sys, math       # load system and math module\n', 'r = float(sys.argv[1]) # extract the 1st command-line arg.\n', 's = math.sin(r)\n', 'print "Hello, World! sin(" + str(r) + ")=" + str(s)\n'],
   'resfile' : <open file 'perl -pe '' hw.py', mode 'r' at 0x402346e0>,
   'root' : '/work/scripting/doc',
   'setcheckinterval' : <built-in function setcheckinterval>,
   'setdlopenflags' : <built-in function setdlopenflags>,
   'setprofile' : <built-in function setprofile>,
   'setrecursionlimit' : <built-in function setrecursionlimit>,
   'settrace' : <built-in function settrace>,
   'shutil' : <module 'shutil' from '/usr/lib/python2.3/shutil.pyc'>,
   'stat' : <module 'stat' from '/usr/lib/python2.3/stat.pyc'>,
   'statistics' : <function statistics at 0x40823684>,
   'stderr' : <open file '<stderr>', mode 'w' at 0x401e40a0>,
   'stdin' : <open file '<stdin>', mode 'r' at 0x401e4020>,
   'stdout' : <open file '<stdout>', mode 'w' at 0x401e4060>,
   'string' : <module 'string' from '/usr/lib/python2.3/string.pyc'>,
   'swap' : <function swap at 0x408236bc>,
   'sys' : <module 'sys' (built-in)>,
   'tail' : 'hw.pl',
   'v1' : 1.3,
   'v2' : 'some text',
   'v3' : 9,
   'value' : '9.8',
   'version' : '2.3.3 (#2, Jan  4 2004, 12:24:16) \n[GCC 3.3.3 20031229 (prerelease) (Debian)]',
   'version_info' : (2, 3, 3, 'final', 0),
   'warnoptions' : [],
   'word' : '  no upwinding',
   'words1' : ['iteration', '12:', 'eps=', '1.245E-05'],
   'words2' : ['.myc_12', 'displacement', 'u(x,3.1415)', '  no upwinding'],
   'write' : <function write at 0x4082387c>,
   },

{
   'a' : 4,
   'b' : {
       'c' : 'some',
       'd' : 77,
       },
   'e' : {
       'f' : {
           'g' : 1,
           'h' : 2,
           },
       'i' : 4,
       },
   },

complex roots: (2-1.41421356237j) (2+1.41421356237j)

regex:

[  just a string   with leading and trailing white space   ]
[just a string   with leading and trailing white space   ]
[just a string   with leading and trailing white space]

comments= []
comments= ['# a comment', '# another comment', '# third comment']
points2= [[ 0.          3.        ]
 [ 0.1         3.57883668]
 [ 0.2         4.03471218]
 [ 0.3         4.26407817]
 [ 0.4         4.19914721]
 [ 0.5         3.81859485]
 [ 0.6         3.15092636]
 [ 0.7         2.2699763 ]
 [ 0.8         1.28325171]
 [ 0.9         0.31495911]
 [ 1.         -0.51360499]
 [ 1.1        -1.10320415]
 [ 1.2        -1.39232922]
 [ 1.3        -1.36690931]
 [ 1.4        -1.06253328]
 [ 1.5        -0.558831  ]
 [ 1.6         0.03309841]
 [ 1.7         0.5882267 ]
 [ 1.8         0.98733573]
 [ 1.9         1.13583934]]
trying urlretrieve: No Internet connection
trying urlopen: No Internet connection
finished
CPU time of commontasks.py: 2.4 seconds on hplx30 i686, Linux


#### Test: ./tests.verify running hw.py 1.2
Hello, World! sin(1.2)=0.932039085967
CPU time of hw.py: 0.1 seconds on hplx30 i686, Linux


#### Test: ./tests.verify running datatrans1.py .datatrans_infile tmp1file
CPU time of datatrans1.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp1file ------
0.1   5.36092e-01
0.2   3.12343e+00
0.3   5.87269e+00
0.4   3.12343e+00

#### Test: ./tests.verify running datatrans2.py .datatrans_infile tmp2file
CPU time of datatrans2.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp2file ------
0.1   5.36092e-01
0.2   3.12343e+00
0.3   5.87269e+00
0.4   3.12343e+00

#### Test: ./tests.verify running datatrans3a.py .datatrans_infile tmp3afile
CPU time of datatrans3a.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp3afile ------
0.1	0.536092209007	
0.2	3.12343489619	
0.3	5.87269405137	
0.4	3.12343489619	

#### Test: ./tests.verify running datatrans3b.py .datatrans_infile tmp3bfile
CPU time of datatrans3b.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp3bfile ------
0.1 0.536092 
0.2 3.12343 
0.3 5.87269 
0.4 3.12343 

#### Test: ./tests.verify running convert1.py .convert_infile1
CPU time of convert1.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp-measurements.dat ------
           0  0.00000e+00
         1.5  1.00000e-01
           3  2.00000e-01


----- appending file tmp-model1.dat ------
           0  1.00000e-01
         1.5  1.00000e-01
           3  2.00000e-01


----- appending file tmp-model2.dat ------
           0  1.00000e+00
         1.5  1.88000e-01
           3  2.50000e-01

#### Test: ./tests.verify running convert2.py .convert_infile1
y dictionary:
{'tmp-model2': [1.0, 0.188, 0.25], 'tmp-model1': [0.10000000000000001, 0.10000000000000001, 0.20000000000000001], 'tmp-measurements': [0.0, 0.10000000000000001, 0.20000000000000001]}
CPU time of convert2.py: 0.1 seconds on hplx30 i686, Linux



----- appending file tmp-measurements.dat ------
           0  0.00000e+00
         1.5  1.00000e-01
           3  2.00000e-01


----- appending file tmp-model1.dat ------
           0  1.00000e-01
         1.5  1.00000e-01
           3  2.00000e-01


----- appending file tmp-model2.dat ------
           0  1.00000e+00
         1.5  1.88000e-01
           3  2.50000e-01

#### Test: ./tests.verify running simviz1.py -A 5.0 -tstop 2 -case tmp4
CPU time of simviz1.py: 0.2 seconds on hplx30 i686, Linux



----- appending file tmp4/tmp4.i ------

        1
        0.7
        5
        y
        5
        6.28319
        0.2
        2
        0.05
        

----- appending file tmp4/tmp4.gnuplot ------

set title 'tmp4: m=1 b=0.7 c=5 f(y)=y A=5 w=6.28319 y0=0.2 dt=0.05';
plot 'sim.dat' title 'y(t)' with lines;

set size ratio 0.3 1.5, 1.0;  
# define the postscript output format:
set term postscript eps monochrome dashed 'Times-Roman' 28;
# output file containing the plot:
set output 'tmp4.ps';
# basic plot command
plot 'sim.dat' title 'y(t)' with lines;
# make a plot in PNG format:
set term png small color;
set output 'tmp4.png';
plot 'sim.dat' title 'y(t)' with lines;


----- appending file tmp4/tmp4.ps (just 30 lines) ------
%!PS-Adobe-2.0 EPSF-2.0
%%Title: tmp4.ps
%%Creator: gnuplot 3.7 patchlevel 3
%%CreationDate: Sun Mar 14 11:56:20 2004
%%DocumentFonts: (atend)
%%BoundingBox: 50 50 590 302
%%Orientation: Portrait
%%EndComments
/gnudict 256 dict def
gnudict begin
/Color false def
/Solid false def
/gnulinewidth 5.000 def
/userlinewidth gnulinewidth def
/vshift -93 def
/dl {10 mul} def
/hpt_ 31.5 def
/vpt_ 31.5 def
/hpt hpt_ def
/vpt vpt_ def
/M {moveto} bind def
/L {lineto} bind def
/R {rmoveto} bind def
/V {rlineto} bind def
/vpt2 vpt 2 mul def
/hpt2 hpt 2 mul def
/Lshow { currentpoint stroke M
  0 vshift R show } def
/Rshow { currentpoint stroke M
  dup stringwidth pop neg vshift R show } def

#### Test: ./tests.verify running loop4simviz2.py c 5 30 2 -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot
MPEG ENCODER STATS (1.5b)
------------------------
TIME STARTED:  Sun Mar 14 11:56:51 2004
MACHINE:  unknown
FIRST FILE:  ./tmp_0000.ppm
LAST FILE:  ./tmp_0012.ppm
PATTERN:  i
GOP_SIZE:  30
SLICES PER FRAME:  1
RANGE:  +/-10
PIXEL SEARCH:  HALF
PSEARCH:  LOGARITHMIC
BSEARCH:  CROSS2
QSCALE:  8 10 25
REFERENCE FRAME:  ORIGINAL


Creating new GOP (closed = T) before frame 0
FRAME 0 (I):  0 seconds  (2882160 bits/s output)
FRAME 1 (I):  0 seconds  (2886240 bits/s output)
FRAME 2 (I):  0 seconds  (2940720 bits/s output)
FRAME 3 (I):  0 seconds  (2907120 bits/s output)
FRAME 4 (I):  0 seconds  (2953200 bits/s output)
FRAME 5 (I):  0 seconds  (3005520 bits/s output)
FRAME 6 (I):  0 seconds  (2977680 bits/s output)
FRAME 7 (I):  0 seconds  (3014640 bits/s output)
FRAME 8 (I):  0 seconds  (3012240 bits/s output)
FRAME 9 (I):  0 seconds  (3011280 bits/s output)
FRAME 10 (I):  0 seconds  (3038400 bits/s output)
FRAME 11 (I):  0 seconds  (3008640 bits/s output)
FRAME 12 (I):  0 seconds  (3065280 bits/s output)


TIME COMPLETED:  Sun Mar 14 11:56:52 2004
Total time:  1 seconds

-------------------------
*****I FRAME SUMMARY*****
-------------------------
  Blocks:     4290     (1288738 bits)     (  300 bpb)
  Frames:       13     (1290104 bits)     (99238 bpf)     (99.9% of total)
  Compression:   20:1     (   1.1747 bpp)
  Seconds:          0     (  45.8824 fps)  (  3876141 pps)  (    15141 mps)
---------------------------------------------
Total Compression:   20:1     (   1.1755 bpp)
Total Frames Per Second:  13.000000 (4290 mps)
CPU Time:  45.882353 fps     (15141 mps)
Total Output Bit Rate (30 fps):  2979230 bits/sec
MPEG file created in :  movie.mpeg


======FRAMES READ:  13
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0000.ppm tmp_c_5/tmp_c_5.ps
tmp_c_5/tmp_c_5.ps transformed via gs to tmp_0000.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0001.ppm tmp_c_7/tmp_c_7.ps
tmp_c_7/tmp_c_7.ps transformed via gs to tmp_0001.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0002.ppm tmp_c_9/tmp_c_9.ps
tmp_c_9/tmp_c_9.ps transformed via gs to tmp_0002.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0003.ppm tmp_c_11/tmp_c_11.ps
tmp_c_11/tmp_c_11.ps transformed via gs to tmp_0003.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0004.ppm tmp_c_13/tmp_c_13.ps
tmp_c_13/tmp_c_13.ps transformed via gs to tmp_0004.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0005.ppm tmp_c_15/tmp_c_15.ps
tmp_c_15/tmp_c_15.ps transformed via gs to tmp_0005.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0006.ppm tmp_c_17/tmp_c_17.ps
tmp_c_17/tmp_c_17.ps transformed via gs to tmp_0006.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0007.ppm tmp_c_19/tmp_c_19.ps
tmp_c_19/tmp_c_19.ps transformed via gs to tmp_0007.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0008.ppm tmp_c_21/tmp_c_21.ps
tmp_c_21/tmp_c_21.ps transformed via gs to tmp_0008.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0009.ppm tmp_c_23/tmp_c_23.ps
tmp_c_23/tmp_c_23.ps transformed via gs to tmp_0009.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0010.ppm tmp_c_25/tmp_c_25.ps
tmp_c_25/tmp_c_25.ps transformed via gs to tmp_0010.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0011.ppm tmp_c_27/tmp_c_27.ps
tmp_c_27/tmp_c_27.ps transformed via gs to tmp_0011.ppm (270 Kb)
gs -q -dBATCH -dNOPAUSE -sDEVICE=ppm  -sOutputFile=tmp_0012.ppm tmp_c_29/tmp_c_29.ps
tmp_c_29/tmp_c_29.ps transformed via gs to tmp_0012.ppm (270 Kb)
mpeg movie in output file movie.mpeg
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 5 -case tmp_c_5
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 7 -case tmp_c_7
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 9 -case tmp_c_9
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 11 -case tmp_c_11
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 13 -case tmp_c_13
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 15 -case tmp_c_15
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 17 -case tmp_c_17
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 19 -case tmp_c_19
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 21 -case tmp_c_21
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 23 -case tmp_c_23
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 25 -case tmp_c_25
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 27 -case tmp_c_27
running python simviz2.py -yaxis -0.7 0.7 -A 5.0 -tstop 2 -case tmp4 -noscreenplot -c 29 -case tmp_c_29
converting PNG files to animated GIF:
convert -delay 50 -loop 1000 tmp_c_5/tmp_c_5.png tmp_c_7/tmp_c_7.png tmp_c_9/tmp_c_9.png tmp_c_11/tmp_c_11.png tmp_c_13/tmp_c_13.png tmp_c_15/tmp_c_15.png tmp_c_17/tmp_c_17.png tmp_c_19/tmp_c_19.png tmp_c_21/tmp_c_21.png tmp_c_23/tmp_c_23.png tmp_c_25/tmp_c_25.png tmp_c_27/tmp_c_27.png tmp_c_29/tmp_c_29.png tmp_c.gif
converting PostScript files to an MPEG movie:
ps2mpeg.py tmp_c_5/tmp_c_5.ps tmp_c_7/tmp_c_7.ps tmp_c_9/tmp_c_9.ps tmp_c_11/tmp_c_11.ps tmp_c_13/tmp_c_13.ps tmp_c_15/tmp_c_15.ps tmp_c_17/tmp_c_17.ps tmp_c_19/tmp_c_19.ps tmp_c_21/tmp_c_21.ps tmp_c_23/tmp_c_23.ps tmp_c_25/tmp_c_25.ps tmp_c_27/tmp_c_27.ps tmp_c_29/tmp_c_29.ps
epsmerge -o tmp_c_runs.ps -x 2 -y 3 -par tmp_c_5/tmp_c_5.ps tmp_c_7/tmp_c_7.ps tmp_c_9/tmp_c_9.ps tmp_c_11/tmp_c_11.ps tmp_c_13/tmp_c_13.ps tmp_c_15/tmp_c_15.ps tmp_c_17/tmp_c_17.ps tmp_c_19/tmp_c_19.ps tmp_c_21/tmp_c_21.ps tmp_c_23/tmp_c_23.ps tmp_c_25/tmp_c_25.ps tmp_c_27/tmp_c_27.ps tmp_c_29/tmp_c_29.ps
CPU time of loop4simviz2.py: 29.5 seconds on hplx30 i686, Linux



----- appending file tmp_c_runs.html ------
<HTML><BODY BGCOLOR="white">
<H1>c=5</H1> <IMG SRC="tmp_c_5/tmp_c_5.png">
<H1>c=7</H1> <IMG SRC="tmp_c_7/tmp_c_7.png">
<H1>c=9</H1> <IMG SRC="tmp_c_9/tmp_c_9.png">
<H1>c=11</H1> <IMG SRC="tmp_c_11/tmp_c_11.png">
<H1>c=13</H1> <IMG SRC="tmp_c_13/tmp_c_13.png">
<H1>c=15</H1> <IMG SRC="tmp_c_15/tmp_c_15.png">
<H1>c=17</H1> <IMG SRC="tmp_c_17/tmp_c_17.png">
<H1>c=19</H1> <IMG SRC="tmp_c_19/tmp_c_19.png">
<H1>c=21</H1> <IMG SRC="tmp_c_21/tmp_c_21.png">
<H1>c=23</H1> <IMG SRC="tmp_c_23/tmp_c_23.png">
<H1>c=25</H1> <IMG SRC="tmp_c_25/tmp_c_25.png">
<H1>c=27</H1> <IMG SRC="tmp_c_27/tmp_c_27.png">
<H1>c=29</H1> <IMG SRC="tmp_c_29/tmp_c_29.png">
<H1>Movie</H1> <IMG SRC="tmp_c.gif">
<H1><A HREF="tmp_c.mpeg">MPEG Movie</A></H1>
</BODY></HTML>

#### Test: ./tests.verify running NumPy_basics.py 
zeros(n, Float): <type 'array'> d [ 0.  0.  0.  0.  0.  0.  0.  0.  0.  0.]
zeros(n) <type 'array'> l [0 0 0 0 0 0 0 0 0 0]
arrayrange(-5, 5, 0.5) <type 'array'> d [-5.  -4.5 -4.  -3.5 -3.  -2.5 -2.  -1.5 -1.  -0.5  0.   0.5  1.   1.5  2. 
       2.5  3.   3.5  4.   4.5  5. ]
y = sin(x/2.0)*3.0: <type 'array'> d [-1.79541643 -2.33421959 -2.72789228 -2.95195784 -2.99248496 -2.84695386
      -2.52441295 -2.04491628 -1.43827662 -0.74221188  0.          0.74221188
       1.43827662  2.04491628  2.52441295  2.84695386  2.99248496  2.95195784
       2.72789228  2.33421959  1.79541643]
pl = [0, 1.2, 4, -9.1, 5, 8]; array(pl, typecode=Float) <type 'array'> [ 0.   1.2  4.  -9.1  5.   8. ]

creating arrays of length 1E+07 ... it may take some time...
fromfunction took 5.39 s and arange&sin took 3.17 s for length 10000000
1.2
[  0.  10.]
[[  0.   1.   2.   3.   4.   5.]
 [  6.   7.   8.   9.  10.  11.]
 [ 12.  13.  14.  15.  16.  17.]
 [ 18.  19.  20.  21.  22.  23.]
 [ 24.  25.  26.  27.  28.  29.]]
[[  6.   8.  10.]
 [ 12.  14.  16.]]
[[  2.   4.]
 [ 20.  22.]]
[[  2.   4.]
 [ 20.  22.]]
a[0,0]=2  a[0,1]=6  a[0,2]=12 
a[1,0]=4  a[1,1]=12  a[1,2]=24 
a.shape = (2,3); a= [[  2.   6.  12.]
 [  4.  12.  24.]]
a.shape = (size(a),); a= [  2.   6.  12.   4.  12.  24.]
b = 3*a - 1; b = clip(b, 0.1, 1.0E+20); c = cos(b) [  5.  17.  35.  11.  35.  71.] [ 0.28366219 -0.27516334 -0.90369221  0.0044257  -0.90369221 -0.30902273]
in-place operations:
multiply(a, 3.0, a); a= [  6.  18.  36.  12.  36.  72.]
subtract(a, 1.0, a); a= [  5.  17.  35.  11.  35.  71.]
divide  (a, 3.0, a); a= [  1.66666667   5.66666667  11.66666667   3.66666667  11.66666667  23.66666667]
add     (a, 1.0, a); a= [  2.66666667   6.66666667  12.66666667   4.66666667  12.66666667  24.66666667]
power   (a, 2.0, a); a= [   7.11111111   44.44444444  160.44444444   21.77777778  160.44444444
       608.44444444]
a[2:4] = -1; a[-1] = a[0]; a= [   7.11111111   44.44444444   -1.           -1.          160.44444444
         7.11111111]
a.shape = (3,2); a[:,0] [   7.11111111   -1.          160.44444444]
a[:,1::2] [[ 44.44444444]
 [ -1.        ]
 [  7.11111111]]
transpose(a):  [[   7.11111111   -1.          160.44444444]
 [  44.44444444   -1.            7.11111111]]
b array entries are of type Float so no casting is necessary
arrayrange(-5, 5, 0.5); variable type=<type 'array'> typecode=d
arrayrange(-5, 5, 1); variable type=<type 'array'> typecode=l
arrayrange(-5.0, 5, 1); variable type=<type 'array'> typecode=d
arrayrange(-5, 5, 0.5, Complex); variable type=<type 'array'> typecode=D
real part of x: [-5.  -4.5 -4.  -3.5 -3.  -2.5 -2.  -1.5 -1.  -0.5  0.   0.5  1.   1.5  2. 
       2.5  3.   3.5  4.   4.5]
imaginary part of x: [ 0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.  0.
       0.]
read from ASCII file: a is <type 'array'> and
   a= [[ 1  2  3  4  5  6  7  8  9 10]
 [11 12 13 14 15 16 17 18 19 20]]
read from binary file: a= [[ 1  2  3  4  5  6  7  8  9 10]
 [11 12 13 14 15 16 17 18 19 20]]


--------- random numbers -------------

random number on (0,1): 0.723068520556
unform random number on (-1,1): -0.874106242503
N(0,1) uniform random number: 1.42433423327
mean of 10000 random uniform random numbers:
on (0,1): 0.496834617839 (should be 0.5)
on (-1,1): -0.0021085279876 (should be 0)
generated 10000 N(0,1) samples with
mean 0.00870529 and st.dev. 0.993361 using RandomArray.normal
probability N(0,1) < 1.5: 0.93


--------- linear algebra -------------

correct solution
correct solution
LinearAlgebra.determinant(A) = 1.19047619048e-05
A*A^-1 =  [[  1.00000000e-00   5.59552404e-14  -1.35003120e-13   8.61533067e-14]
 [ -5.32907052e-15   1.00000000e+00  -1.29007915e-13   8.31557045e-14]
 [ -6.38378239e-15   4.48530102e-14   1.00000000e-00   8.01581024e-14]
 [ -6.35602682e-15   3.93018951e-14  -1.19682042e-13   1.00000000e+00]]
Id =  [[1 0 0 0]
 [0 1 0 0]
 [0 0 1 0]
 [0 0 0 1]]
A*A^-1 - Id =  [[ -2.44249065e-15   5.59552404e-14  -1.35003120e-13   8.61533067e-14]
 [ -5.32907052e-15   4.88498131e-14  -1.29007915e-13   8.31557045e-14]
 [ -6.38378239e-15   4.4853ERROR in ./tests.verify: execution failure arose from the command
  NumPy_basics.py  >> /home/work/scripting/src/py/intro/tests.v

CPU time of NumPy_basics.py: 44.5 seconds on hplx30 i686, Linux


#### Test: ./tests.verify running leastsquares.py 
CPU time of leastsquares.py: 0.3 seconds on hplx30 i686, Linux

